package calc_tb_pkg;

   import uvm_pkg::*;
   `include "uvm_macros.svh"
   `include "calc_rst_trans.sv"
   `include "calc_rst_seqr.sv"
   `include "calc_rst_driver.sv"
   `include "calc_rst_agent.sv"
   `include "calc_out_trans.sv"
   `include "calc_req_trans.sv"
   `include "calc_req_seqr.sv"
   `include "calc_req_driver.sv"
   `include "calc_req_monitor.sv"
   `include "calc_req_agent.sv"
   `include "calc_req_scbd.sv"
   `include "calc_req_env.sv"
   `include "calc_reg.sv"
   `include "calc_reg_model.sv"
   `include "calc_reg_adapter.sv"
   `include "calc_reg_env.sv"
   `include "calc_tb_vseqr.sv"
   `include "calc_tb_env.sv"

   `include "seqlib/calc_seq_reset.sv"
   `include "seqlib/calc_seq_base.sv"
   `include "seqlib/calc_seq_ral_base.sv"
   `include "seqlib/calc_seq_store_fetch.sv"
   `include "seqlib/calc_seq_walking_1s_0s.sv"
   `include "seqlib/calc_seq_arith_cmds.sv"
   `include "seqlib/calc_seq_branch.sv"
   `include "seqlib/calc_seq_overflow.sv"
   `include "seqlib/calc_seq_underflow.sv"
   `include "seqlib/calc_seq_ral.sv"
   `include "seqlib/calc_seq_ordering_rules.sv"

   `include "seqlib/vseq_base.sv"
   `include "seqlib/vseq_store_fetch.sv"
   `include "seqlib/vseq_walking_1s_0s.sv" 
   `include "seqlib/vseq_arith_cmds.sv" 
   `include "seqlib/vseq_branch.sv" 
   `include "seqlib/vseq_overflow.sv" 
   `include "seqlib/vseq_underflow.sv" 
   `include "seqlib/vseq_reset.sv" 
   `include "seqlib/vseq_ral.sv" 
   `include "seqlib/vseq_ordering_rules.sv" 
   
   `include "calc_test.sv"

endpackage : calc_tb_pkg